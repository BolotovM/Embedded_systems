module firstproject
(
	input logic [3:0] A,
	input logic [3:0] B,
	output logic [7:0] C
);
logic [7:0] m;
always_comb
case({A,B})
'b00010001: m <= 1;
'b00010010: m <= 2;
'b00010011: m <= 3;
'b00010100: m <= 4;
'b00010101: m <= 5;
'b00010110: m <= 6;
'b00010111: m <= 7;
'b00011000: m <= 8;
'b00011001: m <= 9;
'b00011010: m <= 10;
'b00011011: m <= 11;
'b00011100: m <= 12;
'b00011101: m <= 13;
'b00011110: m <= 14;
'b00011111: m <= 15;

'b00100001: m <= 2;
'b00100010: m <= 4;
'b00100011: m <= 6;
'b00100100: m <= 8;
'b00100101: m <= 10;
'b00100110: m <= 12;
'b00100111: m <= 14;
'b00101000: m <= 16;
'b00101001: m <= 18;
'b00101010: m <= 20;
'b00101011: m <= 22;
'b00101100: m <= 24;
'b00101101: m <= 26;
'b00101110: m <= 28;
'b00101111: m <= 30;

'b00110001: m <= 3;
'b00110010: m <= 6;
'b00110011: m <= 9;
'b00110100: m <= 12;
'b00110101: m <= 15;
'b00110110: m <= 18;
'b00110111: m <= 21;
'b00111000: m <= 24;
'b00111001: m <= 27;
'b00111010: m <= 30;
'b00111011: m <= 33;
'b00111100: m <= 36;
'b00111101: m <= 39;
'b00111110: m <= 42;
'b00111111: m <= 45;

'b01000001: m <= 4;
'b01000010: m <= 8;
'b01000011: m <= 12;
'b01000100: m <= 16;
'b01000101: m <= 20;
'b01000110: m <= 24;
'b01000111: m <= 28;
'b01001000: m <= 32;
'b01001001: m <= 36;
'b01001010: m <= 40;
'b01001011: m <= 44;
'b01001100: m <= 48;
'b01001101: m <= 52;
'b01001110: m <= 56;
'b01001111: m <= 60;

'b01010001: m <= 5;
'b01010010: m <= 10;
'b01010011: m <= 15;
'b01010100: m <= 20;
'b01010101: m <= 25;
'b01010110: m <= 30;
'b01010111: m <= 35;
'b01011000: m <= 40;
'b01011001: m <= 45;
'b01011010: m <= 50;
'b01011011: m <= 55;
'b01011100: m <= 60;
'b01011101: m <= 65;
'b01011110: m <= 70;
'b01011111: m <= 75;

'b01100001: m <= 6;
'b01100010: m <= 12;
'b01100011: m <= 18;
'b01100100: m <= 24;
'b01100101: m <= 30;
'b01100110: m <= 36;
'b01100111: m <= 42;
'b01101000: m <= 48;
'b01101001: m <= 54;
'b01101010: m <= 60;
'b01101011: m <= 66;
'b01101100: m <= 72;
'b01101101: m <= 78;
'b01101110: m <= 84;
'b01101111: m <= 90;

'b01110001: m <= 7;
'b01110010: m <= 14;
'b01110011: m <= 21;
'b01110100: m <= 28;
'b01110101: m <= 35;
'b01110110: m <= 42;
'b01110111: m <= 49;
'b01111000: m <= 56;
'b01111001: m <= 63;
'b01111010: m <= 70;
'b01111011: m <= 77;
'b01111100: m <= 84;
'b01111101: m <= 91;
'b01111110: m <= 98;
'b01111111: m <= 105;

'b10000001: m <= 8;
'b10000010: m <= 16;
'b10000011: m <= 24;
'b10000100: m <= 32;
'b10000101: m <= 40;
'b10000110: m <= 48;
'b10000111: m <= 56;
'b10001000: m <= 64;
'b10001001: m <= 72;
'b10001010: m <= 80;
'b10001011: m <= 88;
'b10001100: m <= 96;
'b10001101: m <= 104;
'b10001110: m <= 112;
'b10001111: m <= 120;

'b10010001: m <= 9;
'b10010010: m <= 18;
'b10010011: m <= 27;
'b10010100: m <= 36;
'b10010101: m <= 45;
'b10010110: m <= 54;
'b10010111: m <= 63;
'b10011000: m <= 72;
'b10011001: m <= 81;
'b10011010: m <= 90;
'b10011011: m <= 99;
'b10011100: m <= 108;
'b10011101: m <= 117;
'b10011110: m <= 126;
'b10011111: m <= 135;

'b10100001: m <= 10;
'b10100010: m <= 20;
'b10100011: m <= 30;
'b10100100: m <= 40;
'b10100101: m <= 50;
'b10100110: m <= 60;
'b10100111: m <= 70;
'b10101000: m <= 80;
'b10101001: m <= 90;
'b10101010: m <= 100;
'b10101011: m <= 110;
'b10101100: m <= 120;
'b10101101: m <= 130;
'b10101110: m <= 140;
'b10101111: m <= 150;

'b10110001: m <= 11;
'b10110010: m <= 22;
'b10110011: m <= 33;
'b10110100: m <= 44;
'b10110101: m <= 55;
'b10110110: m <= 66;
'b10110111: m <= 77;
'b10111000: m <= 88;
'b10111001: m <= 99;
'b10111010: m <= 110;
'b10111011: m <= 121;
'b10111100: m <= 132;
'b10111101: m <= 143;
'b10111110: m <= 154;
'b10111111: m <= 165;

'b11000001: m <= 12;
'b11000010: m <= 24;
'b11000011: m <= 36;
'b11000100: m <= 48;
'b11000101: m <= 60;
'b11000110: m <= 72;
'b11000111: m <= 84;
'b11001000: m <= 96;
'b11001001: m <= 108;
'b11001010: m <= 120;
'b11001011: m <= 132;
'b11001100: m <= 144;
'b11001101: m <= 156;
'b11001110: m <= 168;
'b11001111: m <= 180;

'b11010001: m <= 13;
'b11010010: m <= 26;
'b11010011: m <= 39;
'b11010100: m <= 52;
'b11010101: m <= 65;
'b11010110: m <= 78;
'b11010111: m <= 91;
'b11011000: m <= 104;
'b11011001: m <= 117;
'b11011010: m <= 130;
'b11011011: m <= 143;
'b11011100: m <= 156;
'b11011101: m <= 169;
'b11011110: m <= 182;
'b11011111: m <= 195;

'b11100001: m <= 14;
'b11100010: m <= 28;
'b11100011: m <= 42;
'b11100100: m <= 56;
'b11100101: m <= 70;
'b11100110: m <= 84;
'b11100111: m <= 98;
'b11101000: m <= 112;
'b11101001: m <= 126;
'b11101010: m <= 140;
'b11101011: m <= 154;
'b11101100: m <= 168;
'b11101101: m <= 182;
'b11101110: m <= 196;
'b11101111: m <= 210;

'b11110001: m <= 15;
'b11110010: m <= 30;
'b11110011: m <= 45;
'b11110100: m <= 60;
'b11110101: m <= 75;
'b11110110: m <= 90;
'b11110111: m <= 105;
'b11111000: m <= 120;
'b11111001: m <= 135;
'b11111010: m <= 150;
'b11111011: m <= 165;
'b11111100: m <= 180;
'b11111101: m <= 195;
'b11111110: m <= 210;
'b11111111: m <= 225;
default: m <= 0;
endcase
assign C = m;
endmodule